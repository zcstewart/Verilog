//Module:		adder
//Input:			[15:0] dataa, [15:0]
//Output:		[15:0] sum

module adder(input [15:0] dataa, datab, output [15:0] sum);
					assign sum = dataa + datab;
endmodule
